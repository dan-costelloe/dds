library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
entity dds is
    Port ( clk : in STD_LOGIC;
           ctrl_word : in STD_LOGIC_VECTOR (7 downto 0);
           data_out : out STD_LOGIC_VECTOR (15 downto 0));
end dds;

architecture Behavioral of dds is
    signal count : unsigned(7 downto 0) := (others=>'0');
    type lut is array (255 downto 0) of integer;
    signal lut_data : unsigned(15 downto 0) := (others=>'0');
    
    constant sine_lut : lut := (
        32768,33575,34382,35187,35992,36794,37594,38391,39185,39975,40760,41540,
        42316,43085,43848,44604,45354,46095,46829,47554,48270,48976,49673,50359,
        51035,51700,52353,52994,53623,54240,54843,55433,56009,56571,57118,57651,
        58169,58671,59158,59628,60083,60520,60941,61345,61731,62100,62451,62784,
        63098,63395,63672,63931,64171,64392,64594,64776,64939,65083,65207,65311,
        65395,65460,65505,65529,65534,65519,65485,65430,65355,65261,65147,65014,
        64860,64688,64495,64284,64054,63804,63536,63249,62943,62619,62277,61918,
        61540,61145,60733,60303,59858,59395,58917,58422,57912,57387,56847,56292,
        55723,55139,54543,53933,53310,52675,52028,51369,50699,50017,49326,48624,
        47913,47192,46463,45725,44980,44227,43467,42701,41929,41151,40368,39580,
        38789,37993,37195,36393,35590,34785,33978,33171,32364,31557,30750,29945,
        29142,28340,27542,26746,25955,25167,24384,23606,22834,22068,21308,20555,
        19810,19072,18343,17622,16911,16209,15518,14836,14166,13507,12860,12225,
        11602,10992,10396,9812,9243,8688,8148,7623,7113,6618,6140,5677,
        5232,4802,4390,3995,3617,3258,2916,2592,2286,1999,1731,1481,
        1251,1040,847,675,521,388,274,180,105,50,16,1,
        6,30,75,140,224,328,452,596,759,941,1143,1364,
        1604,1863,2140,2437,2751,3084,3435,3804,4190,4594,5015,5452,
        5907,6377,6864,7366,7884,8417,8964,9526,10102,10692,11295,11912,
        12541,13182,13835,14500,15176,15862,16559,17265,17981,18706,19440,20181,
        20931,21687,22450,23219,23995,24775,25560,26350,27144,27941,28741,29543,
        30348,31153,31960,32768
    );
begin

COUNTER_8_BIT : process (clk)
begin
    if (clk'event and clk = '1') then
            count <= count + unsigned(ctrl_word);
    end if;
end process;

SINE_LOOKUP : process (clk)
begin
    if (clk'event and clk = '1') then
            data_out <= std_logic_vector(to_unsigned(sine_lut(to_integer(count)),lut_data'length));
    end if;
end process;

				
end Behavioral;
